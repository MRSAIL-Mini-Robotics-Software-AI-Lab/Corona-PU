library IEEE; 
 use IEEE.STD_LOGIC_1164.ALL; 
 use IEEE.numeric_std.ALL; 
 
 entity ROM is 
 port( 
 address : in std_logic_vector(15 downto 0); 
 ROM_tick : in std_logic ; 
 from_ROM: out std_logic_vector(55 downto 0); 
 read_address: in std_logic  
 ); 
 end ROM; 
 
 architecture Behavioral of ROM is 
 -- all data should be declared here as constants as given bellow 
constant data0 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000000000000000000000000" ;
constant data1 : std_logic_vector (55 downto 0) := "00011000010001011000000000000000000000010000000000000001" ;
constant data2 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000000110000000000000011" ;
constant data3 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000001000000000000000100" ;
constant data4 : std_logic_vector (55 downto 0) := "00000011000000000000001100000000000001000000000000000010" ;
constant data5 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000001000000000000000100" ;
constant data6 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000001010000000000000101" ;
constant data7 : std_logic_vector (55 downto 0) := "00000011000000000000010000000000000001010000000000000011" ;
constant data8 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000001010000000000000101" ;
constant data9 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000001100000000000000110" ;
constant data10 : std_logic_vector (55 downto 0) := "00000011000000000000010100000000000001100000000000000100" ;
constant data11 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000001010000000000000101" ;
constant data12 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000001100000000000000110" ;
constant data13 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000001110000000000000111" ;
constant data14 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000010010000000000001001" ;
constant data15 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000010100000000000001010" ;
constant data16 : std_logic_vector (55 downto 0) := "00000011000000000000100100000000000010100000000000001000" ;
constant data17 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000010100000000000001010" ;
constant data18 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000010110000000000001011" ;
constant data19 : std_logic_vector (55 downto 0) := "00000011000000000000101000000000000010110000000000001001" ;
constant data20 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000010100000000000001010" ;
constant data21 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000010110000000000001011" ;
constant data22 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000011000000000000001100" ;
constant data23 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000011010000000000001101" ;
constant data24 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000011110000000000001111" ;
constant data25 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000100000000000000010000" ;
constant data26 : std_logic_vector (55 downto 0) := "00000011000000000000111100000000000100000000000000001110" ;
constant data27 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000011110000000000001111" ;
constant data28 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000100000000000000010000" ;
constant data29 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000100100000000000010010" ;
constant data30 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000100110000000000010011" ;
constant data31 : std_logic_vector (55 downto 0) := "00000011000000000001001000000000000100110000000000010001" ;
constant data32 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000100100000000000010010" ;
constant data33 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000101000000000000010100" ;
constant data34 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000101010000000000010101" ;
constant data35 : std_logic_vector (55 downto 0) := "00000011000000000001010000000000000101010000000000010011" ;
constant data36 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000101000000000000010100" ;
constant data37 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000101010000000000010101" ;
constant data38 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000101110000000000010111" ;
constant data39 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000110000000000000011000" ;
constant data40 : std_logic_vector (55 downto 0) := "00000011000000000001011100000000000110000000000000010110" ;
constant data41 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000110000000000000011000" ;
constant data42 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000110010000000000011001" ;
constant data43 : std_logic_vector (55 downto 0) := "00000011000000000001100000000000000110010000000000010111" ;
constant data44 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000110000000000000011000" ;
constant data45 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000110010000000000011001" ;
constant data46 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000110100000000000011010" ;
constant data47 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000110110000000000011011" ;
constant data48 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000111010000000000011101" ;
constant data49 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000111100000000000011110" ;
constant data50 : std_logic_vector (55 downto 0) := "00000011000000000001110100000000000111100000000000011100" ;
constant data51 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000000111010000000000011101" ;
constant data52 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000111100000000000011110" ;
constant data53 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000000111110000000000011111" ;
constant data54 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001000000000000000100000" ;
constant data55 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001000010000000000100001" ;
constant data56 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001000100000000000100010" ;
constant data57 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001000110000000000100011" ;
constant data58 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001001000000000000100100" ;
constant data59 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001001100000000000100110" ;
constant data60 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001001110000000000100111" ;
constant data61 : std_logic_vector (55 downto 0) := "00000011000000000010011000000000001001110000000000100101" ;
constant data62 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001001100000000000100110" ;
constant data63 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000001001110000000000100111" ;
constant data64 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001010000000000000101000" ;
constant data65 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001010010000000000101001" ;
constant data66 : std_logic_vector (55 downto 0) := "00011000010111100100000000000000001010100000000000101010" ;
constant data67 : std_logic_vector (55 downto 0) := "00011000010111001011000000000000001010110000000000101011" ;
constant data68 : std_logic_vector (55 downto 0) := "00011000010110100100000000000000001011000000000000101100" ;
constant data69 : std_logic_vector (55 downto 0) := "00011000010110001011000000000000001011010000000000101101" ;
constant data70 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001011100000000000101110" ;
constant data71 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001011110000000000101111" ;
constant data72 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001100000000000000110000" ;
constant data73 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001100010000000000110001" ;
constant data74 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001100100000000000110010" ;
constant data75 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001100110000000000110011" ;
constant data76 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001101000000000000110100" ;
constant data77 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001101010000000000110101" ;
constant data78 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001101100000000000110110" ;
constant data79 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001101110000000000110111" ;
constant data80 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001110000000000000111000" ;
constant data81 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001110010000000000111001" ;
constant data82 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001110100000000000111010" ;
constant data83 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001110110000000000111011" ;
constant data84 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001111000000000000111100" ;
constant data85 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001111010000000000111101" ;
constant data86 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001111100000000000111110" ;
constant data87 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000001111110000000000111111" ;
constant data88 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010000000000000001000000" ;
constant data89 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010000010000000001000001" ;
constant data90 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010000100000000001000010" ;
constant data91 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010000110000000001000011" ;
constant data92 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010001000000000001000100" ;
constant data93 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010001010000000001000101" ;
constant data94 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010001100000000001000110" ;
constant data95 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010001110000000001000111" ;
constant data96 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010010000000000001001000" ;
constant data97 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010010010000000001001001" ;
constant data98 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010010100000000001001010" ;
constant data99 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010010110000000001001011" ;
constant data100 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010011000000000001001100" ;
constant data101 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010011010000000001001101" ;
constant data102 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010011100000000001001110" ;
constant data103 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010011110000000001001111" ;
constant data104 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100000000000001010000" ;
constant data105 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data106 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100100000000001010010" ;
constant data107 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100110000000001010011" ;
constant data108 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101000000000001010100" ;
constant data109 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101010000000001010101" ;
constant data110 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data111 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data112 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data113 : std_logic_vector (55 downto 0) := "00011000001001111010111000000000010110010000000001011001" ;
constant data114 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110100000000001011010" ;
constant data115 : std_logic_vector (55 downto 0) := "00011000010110001011000000000000010110110000000001011011" ;
constant data116 : std_logic_vector (55 downto 0) := "00000101000000000101100100000000010110010000000001011100" ;
constant data117 : std_logic_vector (55 downto 0) := "00000101000000000101100100000000010111000000000001011100" ;
constant data118 : std_logic_vector (55 downto 0) := "00000101000000000101100100000000010111000000000001011101" ;
constant data119 : std_logic_vector (55 downto 0) := "00000101000000000101100100000000010111010000000001011101" ;
constant data120 : std_logic_vector (55 downto 0) := "00011000010001100000000000000000010111100000000001011110" ;
constant data121 : std_logic_vector (55 downto 0) := "00000111000000000101110000000000010111100000000001011100" ;
constant data122 : std_logic_vector (55 downto 0) := "00011000010101111000000000000000010111100000000001011110" ;
constant data123 : std_logic_vector (55 downto 0) := "00000111000000000101110100000000010111100000000001011101" ;
constant data124 : std_logic_vector (55 downto 0) := "00000011000000000101100100000000010111000000000001011100" ;
constant data125 : std_logic_vector (55 downto 0) := "00000001000000000101110000000000010111010000000001011101" ;
constant data126 : std_logic_vector (55 downto 0) := "00010111000000000101110100000000001111000000000000111100" ;
constant data127 : std_logic_vector (55 downto 0) := "00011000001111000000000000000000010111000000000001011100" ;
constant data128 : std_logic_vector (55 downto 0) := "00000101000000000101100100000000010110010000000001011101" ;
constant data129 : std_logic_vector (55 downto 0) := "00000101000000000101110100000000010111010000000001011110" ;
constant data130 : std_logic_vector (55 downto 0) := "00011000010001000000000000000000010111110000000001011111" ;
constant data131 : std_logic_vector (55 downto 0) := "00000111000000000101110100000000010111110000000001011101" ;
constant data132 : std_logic_vector (55 downto 0) := "00011000010011100000000000000000010111110000000001011111" ;
constant data133 : std_logic_vector (55 downto 0) := "00000111000000000101111000000000010111110000000001011110" ;
constant data134 : std_logic_vector (55 downto 0) := "00000011000000000101110000000000010111010000000001011101" ;
constant data135 : std_logic_vector (55 downto 0) := "00000001000000000101110100000000010111100000000001011101" ;
constant data136 : std_logic_vector (55 downto 0) := "00010111000000000101111000000000001111010000000000111101" ;
constant data137 : std_logic_vector (55 downto 0) := "00011000001001111010100000000000001111000000000000111100" ;
constant data138 : std_logic_vector (55 downto 0) := "00011000001110111111111000000000001111010000000000111101" ;
constant data139 : std_logic_vector (55 downto 0) := "00000101000000000011110000000000001111010000000000111110" ;
constant data140 : std_logic_vector (55 downto 0) := "00000101000000000011110100000000001111010000000000111111" ;
constant data141 : std_logic_vector (55 downto 0) := "00000101000000000011110000000000001111000000000001000000" ;
constant data142 : std_logic_vector (55 downto 0) := "00000101000000000100000000000000001111000000000001000001" ;
constant data143 : std_logic_vector (55 downto 0) := "00000101000000000100000000000000001111010000000001000010" ;
constant data144 : std_logic_vector (55 downto 0) := "00000101000000000011110000000000001111110000000001000011" ;
constant data145 : std_logic_vector (55 downto 0) := "00000011000000000011111100000000010000010000000001000100" ;
constant data146 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data147 : std_logic_vector (55 downto 0) := "00000011000000000101110000000000001111100000000001000101" ;
constant data148 : std_logic_vector (55 downto 0) := "00000001000000000011111000000000010000100000000001000110" ;
constant data149 : std_logic_vector (55 downto 0) := "00000001000000000011111000000000010000100000000001000111" ;
constant data150 : std_logic_vector (55 downto 0) := "00010111000000000011111100000000010010000000000001001000" ;
constant data151 : std_logic_vector (55 downto 0) := "00000011000000000100000000000000010000110000000001001001" ;
constant data152 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data153 : std_logic_vector (55 downto 0) := "00000011000000000101110000000000001111100000000001001010" ;
constant data154 : std_logic_vector (55 downto 0) := "00010111000000000011110000000000010010110000000001001011" ;
constant data155 : std_logic_vector (55 downto 0) := "00010111000000000011111100000000010011000000000001001100" ;
constant data156 : std_logic_vector (55 downto 0) := "00010110000000000101101000000000100111010000001101111000" ;
constant data157 : std_logic_vector (55 downto 0) := "00000101000000000000001000000000010001000000000000101110" ;
constant data158 : std_logic_vector (55 downto 0) := "00000101000000000000001100000000010001010000000000101111" ;
constant data159 : std_logic_vector (55 downto 0) := "00000101000000000000010000000000010001100000000000110000" ;
constant data160 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data161 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data162 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data163 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data164 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000000101" ;
constant data165 : std_logic_vector (55 downto 0) := "00000101000000000000001000000000010001110000000000101110" ;
constant data166 : std_logic_vector (55 downto 0) := "00000101000000000000001100000000010010000000000000101111" ;
constant data167 : std_logic_vector (55 downto 0) := "00000101000000000000010000000000010010010000000000110000" ;
constant data168 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data169 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data170 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data171 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data172 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000000110" ;
constant data173 : std_logic_vector (55 downto 0) := "00000101000000000000001000000000010010100000000000101110" ;
constant data174 : std_logic_vector (55 downto 0) := "00000101000000000000001100000000010010110000000000101111" ;
constant data175 : std_logic_vector (55 downto 0) := "00000101000000000000010000000000010011000000000000110000" ;
constant data176 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data177 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data178 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000000100000000000000010" ;
constant data179 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000000110000000000000011" ;
constant data180 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000001000000000000000100" ;
constant data181 : std_logic_vector (55 downto 0) := "00000101000000000000011100000000010001000000000000101110" ;
constant data182 : std_logic_vector (55 downto 0) := "00000101000000000000100000000000010001010000000000101111" ;
constant data183 : std_logic_vector (55 downto 0) := "00000101000000000000100100000000010001100000000000110000" ;
constant data184 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data185 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data186 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data187 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data188 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000001010" ;
constant data189 : std_logic_vector (55 downto 0) := "00000101000000000000011100000000010001110000000000101110" ;
constant data190 : std_logic_vector (55 downto 0) := "00000101000000000000100000000000010010000000000000101111" ;
constant data191 : std_logic_vector (55 downto 0) := "00000101000000000000100100000000010010010000000000110000" ;
constant data192 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data193 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data194 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data195 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data196 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000001011" ;
constant data197 : std_logic_vector (55 downto 0) := "00000101000000000000011100000000010010100000000000101110" ;
constant data198 : std_logic_vector (55 downto 0) := "00000101000000000000100000000000010010110000000000101111" ;
constant data199 : std_logic_vector (55 downto 0) := "00000101000000000000100100000000010011000000000000110000" ;
constant data200 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data201 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data202 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000001110000000000000111" ;
constant data203 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000010000000000000001000" ;
constant data204 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000010010000000000001001" ;
constant data205 : std_logic_vector (55 downto 0) := "00000101000000000000110000000000010001000000000000101110" ;
constant data206 : std_logic_vector (55 downto 0) := "00000101000000000000110100000000010001010000000000101111" ;
constant data207 : std_logic_vector (55 downto 0) := "00000101000000000000111000000000010001100000000000110000" ;
constant data208 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data209 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data210 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data211 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data212 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000001111" ;
constant data213 : std_logic_vector (55 downto 0) := "00000101000000000000110000000000010001110000000000101110" ;
constant data214 : std_logic_vector (55 downto 0) := "00000101000000000000110100000000010010000000000000101111" ;
constant data215 : std_logic_vector (55 downto 0) := "00000101000000000000111000000000010010010000000000110000" ;
constant data216 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data217 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data218 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data219 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data220 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000010000" ;
constant data221 : std_logic_vector (55 downto 0) := "00000101000000000000110000000000010010100000000000101110" ;
constant data222 : std_logic_vector (55 downto 0) := "00000101000000000000110100000000010010110000000000101111" ;
constant data223 : std_logic_vector (55 downto 0) := "00000101000000000000111000000000010011000000000000110000" ;
constant data224 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data225 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data226 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000011000000000000001100" ;
constant data227 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000011010000000000001101" ;
constant data228 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000011100000000000001110" ;
constant data229 : std_logic_vector (55 downto 0) := "00000101000000000001000100000000010001000000000000101110" ;
constant data230 : std_logic_vector (55 downto 0) := "00000101000000000001001000000000010001010000000000101111" ;
constant data231 : std_logic_vector (55 downto 0) := "00000101000000000001001100000000010001100000000000110000" ;
constant data232 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data233 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data234 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data235 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data236 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000010100" ;
constant data237 : std_logic_vector (55 downto 0) := "00000101000000000001000100000000010001110000000000101110" ;
constant data238 : std_logic_vector (55 downto 0) := "00000101000000000001001000000000010010000000000000101111" ;
constant data239 : std_logic_vector (55 downto 0) := "00000101000000000001001100000000010010010000000000110000" ;
constant data240 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data241 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data242 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data243 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data244 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000010101" ;
constant data245 : std_logic_vector (55 downto 0) := "00000101000000000001000100000000010010100000000000101110" ;
constant data246 : std_logic_vector (55 downto 0) := "00000101000000000001001000000000010010110000000000101111" ;
constant data247 : std_logic_vector (55 downto 0) := "00000101000000000001001100000000010011000000000000110000" ;
constant data248 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data249 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data250 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000100010000000000010001" ;
constant data251 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000100100000000000010010" ;
constant data252 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000100110000000000010011" ;
constant data253 : std_logic_vector (55 downto 0) := "00000101000000000001011000000000010001000000000000101110" ;
constant data254 : std_logic_vector (55 downto 0) := "00000101000000000001011100000000010001010000000000101111" ;
constant data255 : std_logic_vector (55 downto 0) := "00000101000000000001100000000000010001100000000000110000" ;
constant data256 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data257 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data258 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data259 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data260 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000011001" ;
constant data261 : std_logic_vector (55 downto 0) := "00000101000000000001011000000000010001110000000000101110" ;
constant data262 : std_logic_vector (55 downto 0) := "00000101000000000001011100000000010010000000000000101111" ;
constant data263 : std_logic_vector (55 downto 0) := "00000101000000000001100000000000010010010000000000110000" ;
constant data264 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data265 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data266 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data267 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data268 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000011010" ;
constant data269 : std_logic_vector (55 downto 0) := "00000101000000000001011000000000010010100000000000101110" ;
constant data270 : std_logic_vector (55 downto 0) := "00000101000000000001011100000000010010110000000000101111" ;
constant data271 : std_logic_vector (55 downto 0) := "00000101000000000001100000000000010011000000000000110000" ;
constant data272 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data273 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data274 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000101100000000000010110" ;
constant data275 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000101110000000000010111" ;
constant data276 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000110000000000000011000" ;
constant data277 : std_logic_vector (55 downto 0) := "00000101000000000001101100000000010001000000000000101110" ;
constant data278 : std_logic_vector (55 downto 0) := "00000101000000000001110000000000010001010000000000101111" ;
constant data279 : std_logic_vector (55 downto 0) := "00000101000000000001110100000000010001100000000000110000" ;
constant data280 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data281 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data282 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data283 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data284 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000011110" ;
constant data285 : std_logic_vector (55 downto 0) := "00000101000000000001101100000000010001110000000000101110" ;
constant data286 : std_logic_vector (55 downto 0) := "00000101000000000001110000000000010010000000000000101111" ;
constant data287 : std_logic_vector (55 downto 0) := "00000101000000000001110100000000010010010000000000110000" ;
constant data288 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data289 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data290 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data291 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data292 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000011111" ;
constant data293 : std_logic_vector (55 downto 0) := "00000101000000000001101100000000010010100000000000101110" ;
constant data294 : std_logic_vector (55 downto 0) := "00000101000000000001110000000000010010110000000000101111" ;
constant data295 : std_logic_vector (55 downto 0) := "00000101000000000001110100000000010011000000000000110000" ;
constant data296 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data297 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data298 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000000110110000000000011011" ;
constant data299 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000000111000000000000011100" ;
constant data300 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000000111010000000000011101" ;
constant data301 : std_logic_vector (55 downto 0) := "00000101000000000010000000000000010001000000000000101110" ;
constant data302 : std_logic_vector (55 downto 0) := "00000101000000000010000100000000010001010000000000101111" ;
constant data303 : std_logic_vector (55 downto 0) := "00000101000000000010001000000000010001100000000000110000" ;
constant data304 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data305 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data306 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data307 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data308 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000100011" ;
constant data309 : std_logic_vector (55 downto 0) := "00000101000000000010000000000000010001110000000000101110" ;
constant data310 : std_logic_vector (55 downto 0) := "00000101000000000010000100000000010010000000000000101111" ;
constant data311 : std_logic_vector (55 downto 0) := "00000101000000000010001000000000010010010000000000110000" ;
constant data312 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data313 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data314 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data315 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data316 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000100100" ;
constant data317 : std_logic_vector (55 downto 0) := "00000101000000000010000000000000010010100000000000101110" ;
constant data318 : std_logic_vector (55 downto 0) := "00000101000000000010000100000000010010110000000000101111" ;
constant data319 : std_logic_vector (55 downto 0) := "00000101000000000010001000000000010011000000000000110000" ;
constant data320 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data321 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data322 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000001000000000000000100000" ;
constant data323 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000001000010000000000100001" ;
constant data324 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000001000100000000000100010" ;
constant data325 : std_logic_vector (55 downto 0) := "00000101000000000010010100000000010001000000000000101110" ;
constant data326 : std_logic_vector (55 downto 0) := "00000101000000000010011000000000010001010000000000101111" ;
constant data327 : std_logic_vector (55 downto 0) := "00000101000000000010011100000000010001100000000000110000" ;
constant data328 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110001" ;
constant data329 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001100000000000000110001" ;
constant data330 : std_logic_vector (55 downto 0) := "00010111000000000011000100000000010100100000000001010010" ;
constant data331 : std_logic_vector (55 downto 0) := "00000101000000000011000100000000010110110000000000110001" ;
constant data332 : std_logic_vector (55 downto 0) := "00000001000000000011000100000000001011000000000000101000" ;
constant data333 : std_logic_vector (55 downto 0) := "00000101000000000010010100000000010001110000000000101110" ;
constant data334 : std_logic_vector (55 downto 0) := "00000101000000000010011000000000010010000000000000101111" ;
constant data335 : std_logic_vector (55 downto 0) := "00000101000000000010011100000000010010010000000000110000" ;
constant data336 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000000110010" ;
constant data337 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001100000000000000110010" ;
constant data338 : std_logic_vector (55 downto 0) := "00010111000000000011001000000000010100110000000001010011" ;
constant data339 : std_logic_vector (55 downto 0) := "00000101000000000011001000000000010110110000000000110010" ;
constant data340 : std_logic_vector (55 downto 0) := "00000001000000000011001000000000001011010000000000101001" ;
constant data341 : std_logic_vector (55 downto 0) := "00000101000000000010010100000000010010100000000000101110" ;
constant data342 : std_logic_vector (55 downto 0) := "00000101000000000010011000000000010010110000000000101111" ;
constant data343 : std_logic_vector (55 downto 0) := "00000101000000000010011100000000010011000000000000110000" ;
constant data344 : std_logic_vector (55 downto 0) := "00000001000000000010111000000000001011110000000001010100" ;
constant data345 : std_logic_vector (55 downto 0) := "00000001000000000101010000000000001100000000000001010100" ;
constant data346 : std_logic_vector (55 downto 0) := "00010111000000000101001000000000001001010000000000100101" ;
constant data347 : std_logic_vector (55 downto 0) := "00010111000000000101001100000000001001100000000000100110" ;
constant data348 : std_logic_vector (55 downto 0) := "00010111000000000101010000000000001001110000000000100111" ;
constant data349 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010011010000000001001101" ;
constant data350 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010011100000000001001110" ;
constant data351 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010011110000000001001111" ;
constant data352 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100000000000001010000" ;
constant data353 : std_logic_vector (55 downto 0) := "00010110000000000100110100000001011000100000000101110010" ;
constant data354 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010011100000000001001110" ;
constant data355 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010011110000000001001111" ;
constant data356 : std_logic_vector (55 downto 0) := "00010110000000000100111000000001011001010000000101101110" ;
constant data357 : std_logic_vector (55 downto 0) := "00010100000000000101000000000000000000000000000001010000" ;
constant data358 : std_logic_vector (55 downto 0) := "00010100000000000100111100000000000000000000000001001111" ;
constant data359 : std_logic_vector (55 downto 0) := "00011010000000000101000000000000010011110000000000000000" ;
constant data360 : std_logic_vector (55 downto 0) := "00010101000000000101000000000000000000000000000001010000" ;
constant data361 : std_logic_vector (55 downto 0) := "00010101000000000100111100000000000000000000000001001111" ;
constant data362 : std_logic_vector (55 downto 0) := "00011000001111000000000000000000010111000000000001011100" ;
constant data363 : std_logic_vector (55 downto 0) := "00000001000000000100111100000000010111000000000001001111" ;
constant data364 : std_logic_vector (55 downto 0) := "00001111000000000100111100000000001010100000000001001110" ;
constant data365 : std_logic_vector (55 downto 0) := "00011001000000010110010000000000000000000000000000000000" ;
constant data366 : std_logic_vector (55 downto 0) := "00011000001111000000000000000000010111000000000001011100" ;
constant data367 : std_logic_vector (55 downto 0) := "00000001000000000101000000000000010111000000000001010000" ;
constant data368 : std_logic_vector (55 downto 0) := "00001111000000000101000000000000001010110000000001001101" ;
constant data369 : std_logic_vector (55 downto 0) := "00011001000000010110000100000000000000000000000000000000" ;
constant data370 : std_logic_vector (55 downto 0) := "00010111000000000000010100000000001100110000000000110011" ;
constant data371 : std_logic_vector (55 downto 0) := "00010111000000000000101000000000001101000000000000110100" ;
constant data372 : std_logic_vector (55 downto 0) := "00010111000000000000011000000000001101010000000000110101" ;
constant data373 : std_logic_vector (55 downto 0) := "00010111000000000000101100000000001101100000000000110110" ;
constant data374 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data375 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data376 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data377 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data378 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data379 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data380 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data381 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data382 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001011111110000000110000001" ;
constant data383 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data384 : std_logic_vector (55 downto 0) := "00011001000000011000001000000000000000000000000000000000" ;
constant data385 : std_logic_vector (55 downto 0) := "00011001000000011000001000000000000000000000000000000000" ;
constant data386 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data387 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data388 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001100001010000000110000111" ;
constant data389 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data390 : std_logic_vector (55 downto 0) := "00011001000000011000100000000000000000000000000000000000" ;
constant data391 : std_logic_vector (55 downto 0) := "00011001000000011000100000000000000000000000000000000000" ;
constant data392 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data393 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data394 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data395 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data396 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data397 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data398 : std_logic_vector (55 downto 0) := "00010110000000000101100000000001100011110000000110011101" ;
constant data399 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data400 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data401 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data402 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data403 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data404 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data405 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data406 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data407 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data408 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data409 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data410 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data411 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data412 : std_logic_vector (55 downto 0) := "00011001000000011000111000000000000000000000000000000000" ;
constant data413 : std_logic_vector (55 downto 0) := "00010111000000000000101000000000001100110000000000110011" ;
constant data414 : std_logic_vector (55 downto 0) := "00010111000000000000111100000000001101000000000000110100" ;
constant data415 : std_logic_vector (55 downto 0) := "00010111000000000000101100000000001101010000000000110101" ;
constant data416 : std_logic_vector (55 downto 0) := "00010111000000000001000000000000001101100000000000110110" ;
constant data417 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data418 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data419 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data420 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data421 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data422 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data423 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data424 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data425 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001101010100000000110101100" ;
constant data426 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data427 : std_logic_vector (55 downto 0) := "00011001000000011010110100000000000000000000000000000000" ;
constant data428 : std_logic_vector (55 downto 0) := "00011001000000011010110100000000000000000000000000000000" ;
constant data429 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data430 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data431 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001101100000000000110110010" ;
constant data432 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data433 : std_logic_vector (55 downto 0) := "00011001000000011011001100000000000000000000000000000000" ;
constant data434 : std_logic_vector (55 downto 0) := "00011001000000011011001100000000000000000000000000000000" ;
constant data435 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data436 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data437 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data438 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data439 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data440 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data441 : std_logic_vector (55 downto 0) := "00010110000000000101100000000001101110100000000111001000" ;
constant data442 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data443 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data444 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data445 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data446 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data447 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data448 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data449 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data450 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data451 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data452 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data453 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data454 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data455 : std_logic_vector (55 downto 0) := "00011001000000011011100100000000000000000000000000000000" ;
constant data456 : std_logic_vector (55 downto 0) := "00010111000000000000111100000000001100110000000000110011" ;
constant data457 : std_logic_vector (55 downto 0) := "00010111000000000001010000000000001101000000000000110100" ;
constant data458 : std_logic_vector (55 downto 0) := "00010111000000000001000000000000001101010000000000110101" ;
constant data459 : std_logic_vector (55 downto 0) := "00010111000000000001010100000000001101100000000000110110" ;
constant data460 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data461 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data462 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data463 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data464 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data465 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data466 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data467 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data468 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001110101010000000111010111" ;
constant data469 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data470 : std_logic_vector (55 downto 0) := "00011001000000011101100000000000000000000000000000000000" ;
constant data471 : std_logic_vector (55 downto 0) := "00011001000000011101100000000000000000000000000000000000" ;
constant data472 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data473 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data474 : std_logic_vector (55 downto 0) := "00010110000000000101010100000001110110110000000111011101" ;
constant data475 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data476 : std_logic_vector (55 downto 0) := "00011001000000011101111000000000000000000000000000000000" ;
constant data477 : std_logic_vector (55 downto 0) := "00011001000000011101111000000000000000000000000000000000" ;
constant data478 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data479 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data480 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data481 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data482 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data483 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data484 : std_logic_vector (55 downto 0) := "00010110000000000101100000000001111001010000000111110011" ;
constant data485 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data486 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data487 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data488 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data489 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data490 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data491 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data492 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data493 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data494 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data495 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data496 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data497 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data498 : std_logic_vector (55 downto 0) := "00011001000000011110010000000000000000000000000000000000" ;
constant data499 : std_logic_vector (55 downto 0) := "00010111000000000001010000000000001100110000000000110011" ;
constant data500 : std_logic_vector (55 downto 0) := "00010111000000000000010100000000001101000000000000110100" ;
constant data501 : std_logic_vector (55 downto 0) := "00010111000000000001010100000000001101010000000000110101" ;
constant data502 : std_logic_vector (55 downto 0) := "00010111000000000000011000000000001101100000000000110110" ;
constant data503 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data504 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data505 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data506 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data507 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data508 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data509 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data510 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data511 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010000000000000001000000010" ;
constant data512 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data513 : std_logic_vector (55 downto 0) := "00011001000000100000001100000000000000000000000000000000" ;
constant data514 : std_logic_vector (55 downto 0) := "00011001000000100000001100000000000000000000000000000000" ;
constant data515 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data516 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data517 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010000001100000001000001000" ;
constant data518 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data519 : std_logic_vector (55 downto 0) := "00011001000000100000100100000000000000000000000000000000" ;
constant data520 : std_logic_vector (55 downto 0) := "00011001000000100000100100000000000000000000000000000000" ;
constant data521 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data522 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data523 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data524 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data525 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data526 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data527 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010000100000000001000011110" ;
constant data528 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data529 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data530 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data531 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data532 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data533 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data534 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data535 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data536 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data537 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data538 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data539 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data540 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data541 : std_logic_vector (55 downto 0) := "00011001000000100000111100000000000000000000000000000000" ;
constant data542 : std_logic_vector (55 downto 0) := "00010111000000000001100100000000001100110000000000110011" ;
constant data543 : std_logic_vector (55 downto 0) := "00010111000000000001111000000000001101000000000000110100" ;
constant data544 : std_logic_vector (55 downto 0) := "00010111000000000001101000000000001101010000000000110101" ;
constant data545 : std_logic_vector (55 downto 0) := "00010111000000000001111100000000001101100000000000110110" ;
constant data546 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data547 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data548 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data549 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data550 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data551 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data552 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data553 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data554 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010001010110000001000101101" ;
constant data555 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data556 : std_logic_vector (55 downto 0) := "00011001000000100010111000000000000000000000000000000000" ;
constant data557 : std_logic_vector (55 downto 0) := "00011001000000100010111000000000000000000000000000000000" ;
constant data558 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data559 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data560 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010001100010000001000110011" ;
constant data561 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data562 : std_logic_vector (55 downto 0) := "00011001000000100011010000000000000000000000000000000000" ;
constant data563 : std_logic_vector (55 downto 0) := "00011001000000100011010000000000000000000000000000000000" ;
constant data564 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data565 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data566 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data567 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data568 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data569 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data570 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010001110110000001001001001" ;
constant data571 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data572 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data573 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data574 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data575 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data576 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data577 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data578 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data579 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data580 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data581 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data582 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data583 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data584 : std_logic_vector (55 downto 0) := "00011001000000100011101000000000000000000000000000000000" ;
constant data585 : std_logic_vector (55 downto 0) := "00010111000000000001111000000000001100110000000000110011" ;
constant data586 : std_logic_vector (55 downto 0) := "00010111000000000010001100000000001101000000000000110100" ;
constant data587 : std_logic_vector (55 downto 0) := "00010111000000000001111100000000001101010000000000110101" ;
constant data588 : std_logic_vector (55 downto 0) := "00010111000000000010010000000000001101100000000000110110" ;
constant data589 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data590 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data591 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data592 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data593 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data594 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data595 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data596 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data597 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010010101100000001001011000" ;
constant data598 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data599 : std_logic_vector (55 downto 0) := "00011001000000100101100100000000000000000000000000000000" ;
constant data600 : std_logic_vector (55 downto 0) := "00011001000000100101100100000000000000000000000000000000" ;
constant data601 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data602 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data603 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010010111000000001001011110" ;
constant data604 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data605 : std_logic_vector (55 downto 0) := "00011001000000100101111100000000000000000000000000000000" ;
constant data606 : std_logic_vector (55 downto 0) := "00011001000000100101111100000000000000000000000000000000" ;
constant data607 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data608 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data609 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data610 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data611 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data612 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data613 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010011001100000001001110100" ;
constant data614 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data615 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data616 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data617 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data618 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data619 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data620 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data621 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data622 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data623 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data624 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data625 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data626 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data627 : std_logic_vector (55 downto 0) := "00011001000000100110010100000000000000000000000000000000" ;
constant data628 : std_logic_vector (55 downto 0) := "00010111000000000010001100000000001100110000000000110011" ;
constant data629 : std_logic_vector (55 downto 0) := "00010111000000000010100000000000001101000000000000110100" ;
constant data630 : std_logic_vector (55 downto 0) := "00010111000000000010010000000000001101010000000000110101" ;
constant data631 : std_logic_vector (55 downto 0) := "00010111000000000010100100000000001101100000000000110110" ;
constant data632 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data633 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data634 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data635 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data636 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data637 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data638 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data639 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data640 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010100000010000001010000011" ;
constant data641 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data642 : std_logic_vector (55 downto 0) := "00011001000000101000010000000000000000000000000000000000" ;
constant data643 : std_logic_vector (55 downto 0) := "00011001000000101000010000000000000000000000000000000000" ;
constant data644 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data645 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data646 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010100001110000001010001001" ;
constant data647 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data648 : std_logic_vector (55 downto 0) := "00011001000000101000101000000000000000000000000000000000" ;
constant data649 : std_logic_vector (55 downto 0) := "00011001000000101000101000000000000000000000000000000000" ;
constant data650 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data651 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data652 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data653 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data654 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data655 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data656 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010100100010000001010011111" ;
constant data657 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data658 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data659 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data660 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data661 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data662 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data663 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data664 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data665 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data666 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data667 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data668 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data669 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data670 : std_logic_vector (55 downto 0) := "00011001000000101001000000000000000000000000000000000000" ;
constant data671 : std_logic_vector (55 downto 0) := "00010111000000000010100000000000001100110000000000110011" ;
constant data672 : std_logic_vector (55 downto 0) := "00010111000000000001100100000000001101000000000000110100" ;
constant data673 : std_logic_vector (55 downto 0) := "00010111000000000010100100000000001101010000000000110101" ;
constant data674 : std_logic_vector (55 downto 0) := "00010111000000000001101000000000001101100000000000110110" ;
constant data675 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data676 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data677 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data678 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data679 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data680 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data681 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data682 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data683 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010101011000000001010101110" ;
constant data684 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data685 : std_logic_vector (55 downto 0) := "00011001000000101010111100000000000000000000000000000000" ;
constant data686 : std_logic_vector (55 downto 0) := "00011001000000101010111100000000000000000000000000000000" ;
constant data687 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data688 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data689 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010101100100000001010110100" ;
constant data690 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data691 : std_logic_vector (55 downto 0) := "00011001000000101011010100000000000000000000000000000000" ;
constant data692 : std_logic_vector (55 downto 0) := "00011001000000101011010100000000000000000000000000000000" ;
constant data693 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data694 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data695 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data696 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data697 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data698 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data699 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010101111000000001011001010" ;
constant data700 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data701 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data702 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data703 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data704 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data705 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data706 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data707 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data708 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data709 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data710 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data711 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data712 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data713 : std_logic_vector (55 downto 0) := "00011001000000101011101100000000000000000000000000000000" ;
constant data714 : std_logic_vector (55 downto 0) := "00010111000000000000010100000000001100110000000000110011" ;
constant data715 : std_logic_vector (55 downto 0) := "00010111000000000001100100000000001101000000000000110100" ;
constant data716 : std_logic_vector (55 downto 0) := "00010111000000000000011000000000001101010000000000110101" ;
constant data717 : std_logic_vector (55 downto 0) := "00010111000000000001101000000000001101100000000000110110" ;
constant data718 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data719 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data720 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data721 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data722 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data723 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data724 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data725 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data726 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010110101110000001011011001" ;
constant data727 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data728 : std_logic_vector (55 downto 0) := "00011001000000101101101000000000000000000000000000000000" ;
constant data729 : std_logic_vector (55 downto 0) := "00011001000000101101101000000000000000000000000000000000" ;
constant data730 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data731 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data732 : std_logic_vector (55 downto 0) := "00010110000000000101010100000010110111010000001011011111" ;
constant data733 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data734 : std_logic_vector (55 downto 0) := "00011001000000101110000000000000000000000000000000000000" ;
constant data735 : std_logic_vector (55 downto 0) := "00011001000000101110000000000000000000000000000000000000" ;
constant data736 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data737 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data738 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data739 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data740 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data741 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data742 : std_logic_vector (55 downto 0) := "00010110000000000101100000000010111001110000001011110101" ;
constant data743 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data744 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data745 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data746 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data747 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data748 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data749 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data750 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data751 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data752 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data753 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data754 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data755 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data756 : std_logic_vector (55 downto 0) := "00011001000000101110011000000000000000000000000000000000" ;
constant data757 : std_logic_vector (55 downto 0) := "00010111000000000000101000000000001100110000000000110011" ;
constant data758 : std_logic_vector (55 downto 0) := "00010111000000000001111000000000001101000000000000110100" ;
constant data759 : std_logic_vector (55 downto 0) := "00010111000000000000101100000000001101010000000000110101" ;
constant data760 : std_logic_vector (55 downto 0) := "00010111000000000001111100000000001101100000000000110110" ;
constant data761 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data762 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data763 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data764 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data765 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data766 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data767 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data768 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data769 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011000000100000001100000100" ;
constant data770 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data771 : std_logic_vector (55 downto 0) := "00011001000000110000010100000000000000000000000000000000" ;
constant data772 : std_logic_vector (55 downto 0) := "00011001000000110000010100000000000000000000000000000000" ;
constant data773 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data774 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data775 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011000010000000001100001010" ;
constant data776 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data777 : std_logic_vector (55 downto 0) := "00011001000000110000101100000000000000000000000000000000" ;
constant data778 : std_logic_vector (55 downto 0) := "00011001000000110000101100000000000000000000000000000000" ;
constant data779 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data780 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data781 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data782 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data783 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data784 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data785 : std_logic_vector (55 downto 0) := "00010110000000000101100000000011000100100000001100100000" ;
constant data786 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data787 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data788 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data789 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data790 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data791 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data792 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data793 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data794 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data795 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data796 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data797 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data798 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data799 : std_logic_vector (55 downto 0) := "00011001000000110001000100000000000000000000000000000000" ;
constant data800 : std_logic_vector (55 downto 0) := "00010111000000000000111100000000001100110000000000110011" ;
constant data801 : std_logic_vector (55 downto 0) := "00010111000000000010001100000000001101000000000000110100" ;
constant data802 : std_logic_vector (55 downto 0) := "00010111000000000001000000000000001101010000000000110101" ;
constant data803 : std_logic_vector (55 downto 0) := "00010111000000000010010000000000001101100000000000110110" ;
constant data804 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data805 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data806 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data807 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data808 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data809 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data810 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data811 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data812 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011001011010000001100101111" ;
constant data813 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data814 : std_logic_vector (55 downto 0) := "00011001000000110011000000000000000000000000000000000000" ;
constant data815 : std_logic_vector (55 downto 0) := "00011001000000110011000000000000000000000000000000000000" ;
constant data816 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data817 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data818 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011001100110000001100110101" ;
constant data819 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data820 : std_logic_vector (55 downto 0) := "00011001000000110011011000000000000000000000000000000000" ;
constant data821 : std_logic_vector (55 downto 0) := "00011001000000110011011000000000000000000000000000000000" ;
constant data822 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data823 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data824 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data825 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data826 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data827 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data828 : std_logic_vector (55 downto 0) := "00010110000000000101100000000011001111010000001101001011" ;
constant data829 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data830 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data831 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data832 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data833 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data834 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data835 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data836 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data837 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data838 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data839 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data840 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data841 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data842 : std_logic_vector (55 downto 0) := "00011001000000110011110000000000000000000000000000000000" ;
constant data843 : std_logic_vector (55 downto 0) := "00010111000000000001010000000000001100110000000000110011" ;
constant data844 : std_logic_vector (55 downto 0) := "00010111000000000010100000000000001101000000000000110100" ;
constant data845 : std_logic_vector (55 downto 0) := "00010111000000000001010100000000001101010000000000110101" ;
constant data846 : std_logic_vector (55 downto 0) := "00010111000000000010100100000000001101100000000000110110" ;
constant data847 : std_logic_vector (55 downto 0) := "00000011000000000011010000000000001100110000000000110111" ;
constant data848 : std_logic_vector (55 downto 0) := "00000011000000000011011000000000001101010000000000111000" ;
constant data849 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data850 : std_logic_vector (55 downto 0) := "00000111000000000011011100000000010111000000000000110111" ;
constant data851 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data852 : std_logic_vector (55 downto 0) := "00000111000000000011100000000000010111000000000000111000" ;
constant data853 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data854 : std_logic_vector (55 downto 0) := "00001101000000000011011100000000010111000000000001010101" ;
constant data855 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011010110000000001101011010" ;
constant data856 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001101110000000000110111" ;
constant data857 : std_logic_vector (55 downto 0) := "00011001000000110101101100000000000000000000000000000000" ;
constant data858 : std_logic_vector (55 downto 0) := "00011001000000110101101100000000000000000000000000000000" ;
constant data859 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010111000000000001011100" ;
constant data860 : std_logic_vector (55 downto 0) := "00001101000000000011100000000000010111000000000001010101" ;
constant data861 : std_logic_vector (55 downto 0) := "00010110000000000101010100000011010111100000001101100000" ;
constant data862 : std_logic_vector (55 downto 0) := "00011000000101000001100100000000001110000000000000111000" ;
constant data863 : std_logic_vector (55 downto 0) := "00011001000000110110000100000000000000000000000000000000" ;
constant data864 : std_logic_vector (55 downto 0) := "00011001000000110110000100000000000000000000000000000000" ;
constant data865 : std_logic_vector (55 downto 0) := "00010111000000000011001100000000001110100000000000111010" ;
constant data866 : std_logic_vector (55 downto 0) := "00010111000000000011010100000000001110110000000000111011" ;
constant data867 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010100010000000001010001" ;
constant data868 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101110000000001010111" ;
constant data869 : std_logic_vector (55 downto 0) := "00011000000000000000000000000000010101100000000001010110" ;
constant data870 : std_logic_vector (55 downto 0) := "00011000000000000000000100000000010110000000000001011000" ;
constant data871 : std_logic_vector (55 downto 0) := "00010110000000000101100000000011011010000000001101110110" ;
constant data872 : std_logic_vector (55 downto 0) := "00000101000000000011100000000000010100010000000001010111" ;
constant data873 : std_logic_vector (55 downto 0) := "00000001000000000101011100000000001110110000000001010111" ;
constant data874 : std_logic_vector (55 downto 0) := "00000101000000000011011100000000010100010000000001010110" ;
constant data875 : std_logic_vector (55 downto 0) := "00000001000000000101011000000000001110100000000001010110" ;
constant data876 : std_logic_vector (55 downto 0) := "00010100000000000101011100000000000000000000000001010111" ;
constant data877 : std_logic_vector (55 downto 0) := "00010100000000000101011000000000000000000000000001010110" ;
constant data878 : std_logic_vector (55 downto 0) := "00011010000000000101011100000000010101100000000000000001" ;
constant data879 : std_logic_vector (55 downto 0) := "00010101000000000101011100000000000000000000000001010111" ;
constant data880 : std_logic_vector (55 downto 0) := "00010101000000000101011000000000000000000000000001010110" ;
constant data881 : std_logic_vector (55 downto 0) := "00011000001110000000000000000000010111000000000001011100" ;
constant data882 : std_logic_vector (55 downto 0) := "00000001000000000101000100000000010111000000000001010001" ;
constant data883 : std_logic_vector (55 downto 0) := "00011000010101100100000000000000010111000000000001011100" ;
constant data884 : std_logic_vector (55 downto 0) := "00001111000000000101000100000000010111000000000001011000" ;
constant data885 : std_logic_vector (55 downto 0) := "00011001000000110110011100000000000000000000000000000000" ;
constant data886 : std_logic_vector (55 downto 0) := "00011011000000000000000000000000000000000000000000000000" ;
constant data887 : std_logic_vector (55 downto 0) := "00011001000000001001110000000000000000000000000000000000" ;
type rom_t is array (natural range <> ) of std_logic_vector  (55 downto 0) ;

constant myrom : rom_t := ( data0,data1,data2,data3,data4,data5,data6,data7,data8,data9,data10,data11,data12,data13,data14,data15,data16,data17,data18,data19,data20,data21,data22,data23,data24,data25,data26,data27,data28,data29,data30,data31,data32,data33,data34,data35,data36,data37,data38,data39,data40,data41,data42,data43,data44,data45,data46,data47,data48,data49,data50,data51,data52,data53,data54,data55,data56,data57,data58,data59,data60,data61,data62,data63,data64,data65,data66,data67,data68,data69,data70,data71,data72,data73,data74,data75,data76,data77,data78,data79,data80,data81,data82,data83,data84,data85,data86,data87,data88,data89,data90,data91,data92,data93,data94,data95,data96,data97,data98,data99,data100,data101,data102,data103,data104,data105,data106,data107,data108,data109,data110,data111,data112,data113,data114,data115,data116,data117,data118,data119,data120,data121,data122,data123,data124,data125,data126,data127,data128,data129,data130,data131,data132,data133,data134,data135,data136,data137,data138,data139,data140,data141,data142,data143,data144,data145,data146,data147,data148,data149,data150,data151,data152,data153,data154,data155,data156,data157,data158,data159,data160,data161,data162,data163,data164,data165,data166,data167,data168,data169,data170,data171,data172,data173,data174,data175,data176,data177,data178,data179,data180,data181,data182,data183,data184,data185,data186,data187,data188,data189,data190,data191,data192,data193,data194,data195,data196,data197,data198,data199,data200,data201,data202,data203,data204,data205,data206,data207,data208,data209,data210,data211,data212,data213,data214,data215,data216,data217,data218,data219,data220,data221,data222,data223,data224,data225,data226,data227,data228,data229,data230,data231,data232,data233,data234,data235,data236,data237,data238,data239,data240,data241,data242,data243,data244,data245,data246,data247,data248,data249,data250,data251,data252,data253,data254,data255,data256,data257,data258,data259,data260,data261,data262,data263,data264,data265,data266,data267,data268,data269,data270,data271,data272,data273,data274,data275,data276,data277,data278,data279,data280,data281,data282,data283,data284,data285,data286,data287,data288,data289,data290,data291,data292,data293,data294,data295,data296,data297,data298,data299,data300,data301,data302,data303,data304,data305,data306,data307,data308,data309,data310,data311,data312,data313,data314,data315,data316,data317,data318,data319,data320,data321,data322,data323,data324,data325,data326,data327,data328,data329,data330,data331,data332,data333,data334,data335,data336,data337,data338,data339,data340,data341,data342,data343,data344,data345,data346,data347,data348,data349,data350,data351,data352,data353,data354,data355,data356,data357,data358,data359,data360,data361,data362,data363,data364,data365,data366,data367,data368,data369,data370,data371,data372,data373,data374,data375,data376,data377,data378,data379,data380,data381,data382,data383,data384,data385,data386,data387,data388,data389,data390,data391,data392,data393,data394,data395,data396,data397,data398,data399,data400,data401,data402,data403,data404,data405,data406,data407,data408,data409,data410,data411,data412,data413,data414,data415,data416,data417,data418,data419,data420,data421,data422,data423,data424,data425,data426,data427,data428,data429,data430,data431,data432,data433,data434,data435,data436,data437,data438,data439,data440,data441,data442,data443,data444,data445,data446,data447,data448,data449,data450,data451,data452,data453,data454,data455,data456,data457,data458,data459,data460,data461,data462,data463,data464,data465,data466,data467,data468,data469,data470,data471,data472,data473,data474,data475,data476,data477,data478,data479,data480,data481,data482,data483,data484,data485,data486,data487,data488,data489,data490,data491,data492,data493,data494,data495,data496,data497,data498,data499,data500,data501,data502,data503,data504,data505,data506,data507,data508,data509,data510,data511,data512,data513,data514,data515,data516,data517,data518,data519,data520,data521,data522,data523,data524,data525,data526,data527,data528,data529,data530,data531,data532,data533,data534,data535,data536,data537,data538,data539,data540,data541,data542,data543,data544,data545,data546,data547,data548,data549,data550,data551,data552,data553,data554,data555,data556,data557,data558,data559,data560,data561,data562,data563,data564,data565,data566,data567,data568,data569,data570,data571,data572,data573,data574,data575,data576,data577,data578,data579,data580,data581,data582,data583,data584,data585,data586,data587,data588,data589,data590,data591,data592,data593,data594,data595,data596,data597,data598,data599,data600,data601,data602,data603,data604,data605,data606,data607,data608,data609,data610,data611,data612,data613,data614,data615,data616,data617,data618,data619,data620,data621,data622,data623,data624,data625,data626,data627,data628,data629,data630,data631,data632,data633,data634,data635,data636,data637,data638,data639,data640,data641,data642,data643,data644,data645,data646,data647,data648,data649,data650,data651,data652,data653,data654,data655,data656,data657,data658,data659,data660,data661,data662,data663,data664,data665,data666,data667,data668,data669,data670,data671,data672,data673,data674,data675,data676,data677,data678,data679,data680,data681,data682,data683,data684,data685,data686,data687,data688,data689,data690,data691,data692,data693,data694,data695,data696,data697,data698,data699,data700,data701,data702,data703,data704,data705,data706,data707,data708,data709,data710,data711,data712,data713,data714,data715,data716,data717,data718,data719,data720,data721,data722,data723,data724,data725,data726,data727,data728,data729,data730,data731,data732,data733,data734,data735,data736,data737,data738,data739,data740,data741,data742,data743,data744,data745,data746,data747,data748,data749,data750,data751,data752,data753,data754,data755,data756,data757,data758,data759,data760,data761,data762,data763,data764,data765,data766,data767,data768,data769,data770,data771,data772,data773,data774,data775,data776,data777,data778,data779,data780,data781,data782,data783,data784,data785,data786,data787,data788,data789,data790,data791,data792,data793,data794,data795,data796,data797,data798,data799,data800,data801,data802,data803,data804,data805,data806,data807,data808,data809,data810,data811,data812,data813,data814,data815,data816,data817,data818,data819,data820,data821,data822,data823,data824,data825,data826,data827,data828,data829,data830,data831,data832,data833,data834,data835,data836,data837,data838,data839,data840,data841,data842,data843,data844,data845,data846,data847,data848,data849,data850,data851,data852,data853,data854,data855,data856,data857,data858,data859,data860,data861,data862,data863,data864,data865,data866,data867,data868,data869,data870,data871,data872,data873,data874,data875,data876,data877,data878,data879,data880,data881,data882,data883,data884,data885,data886,data887);
signal s_ad:integer range 0 to 888 ; 
signal count : integer range 0 to 887 ;
 begin 
 process (ROM_tick) 
 begin 
 if (ROM_tick = '1') then 
 if (read_address = '1') then  
 count <= to_integer(unsigned(address)); 
 elsif ( count < 887 ) then 
 count <= count + 1;  
 end if;  
 end if ; 
 end process ; 
 s_ad <= count; 
 from_ROM <= myrom(s_ad); 
 end Behavioral;